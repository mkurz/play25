hello=Hejsan